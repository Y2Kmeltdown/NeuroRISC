module writeback(

);

endmodule 